// Copyright 2017 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the “License”); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

  logic [31:0]     data_mem[];  // this variable holds the whole memory content
  logic [31:0]     instr_mem[]; // this variable holds the whole memory content
  event            event_mem_load;


`define mem_preload_netlist    //  preloads netlist extraceted memory generated by Vivado
//`define mem_preload_behav      // preloads the behaivioral memories of the PULPino core

`ifdef mem_preload_behav
`undef  mem_preload_netlist
`endif

`ifdef mem_preload_netlist
`undef  mem_preload_behav
`endif

`ifdef mem_preload_behav
  task mem_preload;
    integer      addr;
    integer      mem_addr_dmem;
    integer      mem_addr_pmem;
    integer      mem_addr;
    integer      bidx;
    integer      instr_size;
    integer      instr_width;
    integer      data_size;
    integer      data_width;
    logic [31:0] data_dmem;
    logic [31:0] data_pmem;
    logic [31:0] data;
    string       l2_imem_file;
    string       l2_dmem_file;
    begin
      $display("Preloading memory");

      instr_size   = tb.top_i.core_region_i.instr_mem.mem_gen.sp_ram_wrap_i.RAM_SIZE;
      instr_width = tb.top_i.core_region_i.instr_mem.mem_gen.sp_ram_wrap_i.DATA_WIDTH;

      data_size   = tb.top_i.core_region_i.mem_gen.data_mem.RAM_SIZE;
      data_width = tb.top_i.core_region_i.mem_gen.data_mem.DATA_WIDTH;

      instr_mem = new [instr_size/4];
      data_mem  = new [data_size/4];

      if(!$value$plusargs("l2_imem=%s", l2_imem_file))
         l2_imem_file = "slm_files/l2_stim.slm";

      $display("Preloading instruction memory from %0s", l2_imem_file);
      $readmemh(l2_imem_file, instr_mem);

      if(!$value$plusargs("l2_dmem=%s", l2_dmem_file))
         l2_dmem_file = "slm_files/tcdm_bank0.slm";

      $display("Preloading data memory from %0s", l2_dmem_file);
      $readmemh(l2_dmem_file, data_mem);


      `ifdef mem_preload_behav
        // preload data memory
        for(addr = 0; addr < data_size/4; addr = addr) begin
          for(bidx = 0; bidx < data_width/8; bidx++) begin
            mem_addr = addr / (data_width/32);
            data = data_mem[addr];
            if (bidx%4 == 0)
              tb.top_i.core_region_i.mem_gen.data_mem.sp_ram_i.mem[mem_addr][bidx] = data[ 7: 0];
            else if (bidx%4 == 1)
              tb.top_i.core_region_i.mem_gen.data_mem.sp_ram_i.mem[mem_addr][bidx] = data[15: 8];
            else if (bidx%4 == 2)
              tb.top_i.core_region_i.mem_gen.data_mem.sp_ram_i.mem[mem_addr][bidx] = data[23:16];
            else if (bidx%4 == 3)
              tb.top_i.core_region_i.mem_gen.data_mem.sp_ram_i.mem[mem_addr][bidx] = data[31:24];

            if (bidx%4 == 3) addr++;
          end
        end

        // preload instruction memory
        for(addr = 0; addr < instr_size/4; addr = addr) begin
          for(bidx = 0; bidx < instr_width/8; bidx++) begin
            mem_addr = addr / (instr_width/32);
            data = instr_mem[addr];
            if (bidx%4 == 0)
              tb.top_i.core_region_i.instr_mem.mem_gen.sp_ram_wrap_i.sp_ram_i.mem[mem_addr][bidx] = data[ 7: 0];
            else if (bidx%4 == 1)
              tb.top_i.core_region_i.instr_mem.mem_gen.sp_ram_wrap_i.sp_ram_i.mem[mem_addr][bidx] = data[15: 8];
            else if (bidx%4 == 2)
              tb.top_i.core_region_i.instr_mem.mem_gen.sp_ram_wrap_i.sp_ram_i.mem[mem_addr][bidx] = data[23:16];
            else if (bidx%4 == 3)
              tb.top_i.core_region_i.instr_mem.mem_gen.sp_ram_wrap_i.sp_ram_i.mem[mem_addr][bidx] = data[31:24];

            if (bidx%4 == 3) addr++;
          end
        end
      `endif

    end
  endtask
`endif

`ifdef mem_preload_netlist
  task mem_preload;
    integer      addr;
    integer      mem_addr_dmem;
    integer      mem_addr_pmem;
    integer      mem_addr;
    integer      bidx;
    integer      instr_size;
    integer      instr_width;
    integer      data_size;
    integer      data_width;
    logic [31:0] data_dmem;
    logic [31:0] data_pmem;
    logic [31:0] data;
    string       l2_imem_file;
    string       l2_dmem_file;
    begin
      $display("Preloading memory");

      instr_size = 32768;
      instr_width = 32;

      data_size = 32768;
      data_width = 32;

      instr_mem = new [instr_size/4];
      data_mem  = new [data_size/4];

      if(!$value$plusargs("l2_imem=%s", l2_imem_file))
         l2_imem_file = "slm_files/l2_stim.slm";

      $display("Preloading instruction memory from %0s", l2_imem_file);
      $readmemh(l2_imem_file, instr_mem);

      if(!$value$plusargs("l2_dmem=%s", l2_dmem_file))
         l2_dmem_file = "slm_files/tcdm_bank0.slm";

      $display("Preloading data memory from %0s", l2_dmem_file);
      $readmemh(l2_dmem_file, data_mem);


      // preload data memory
      // preload instruction memory

      `ifdef mem_preload_netlist
        for(addr = 0; addr < data_size/4; addr++) begin
		  #10
          mem_addr_dmem = addr / (data_width/32);
          data_dmem = data_mem[addr];
          force tb.top_i.core_region_i.mem_gen_net.data_mem.addr_i_IBUF = mem_addr_dmem;
          force tb.top_i.core_region_i.mem_gen_net.data_mem.en_i_IBUF   = 1'b1;
          force tb.top_i.core_region_i.mem_gen_net.data_mem.sp_ram_i_i_1_n_0 = 1'b1;
          force tb.top_i.core_region_i.mem_gen_net.data_mem.sp_ram_i_i_2_n_0 = 1'b1;
          force tb.top_i.core_region_i.mem_gen_net.data_mem.sp_ram_i_i_3_n_0 = 1'b1;
          force tb.top_i.core_region_i.mem_gen_net.data_mem.sp_ram_i_i_4_n_0 = 1'b1;
          force tb.top_i.core_region_i.mem_gen_net.data_mem.wdata_i_IBUF = data_dmem;
          mem_addr_pmem = addr / (instr_width/32);
          data_pmem = instr_mem[addr];
          force tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.addr_i_IBUF = mem_addr_pmem;
          force tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.en_i_IBUF   = 1'b1;
          force tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.sp_ram_i_i_1_n_0 = 1'b1;
          force tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.sp_ram_i_i_2_n_0 = 1'b1;
          force tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.sp_ram_i_i_3_n_0 = 1'b1;
          force tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.sp_ram_i_i_4_n_0 = 1'b1;
          force tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.wdata_i_IBUF = data_pmem;
        end
        release tb.top_i.core_region_i.mem_gen_net.data_mem.addr_i_IBUF;
        release tb.top_i.core_region_i.mem_gen_net.data_mem.sp_ram_i_i_1_n_0;
        release tb.top_i.core_region_i.mem_gen_net.data_mem.sp_ram_i_i_2_n_0;
        release tb.top_i.core_region_i.mem_gen_net.data_mem.sp_ram_i_i_3_n_0;
        release tb.top_i.core_region_i.mem_gen_net.data_mem.sp_ram_i_i_4_n_0;
        release tb.top_i.core_region_i.mem_gen_net.data_mem.wdata_i_IBUF;
        release tb.top_i.core_region_i.mem_gen_net.data_mem.en_i_IBUF;

        release tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.addr_i_IBUF;
        release tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.sp_ram_i_i_1_n_0;
        release tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.sp_ram_i_i_2_n_0;
        release tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.sp_ram_i_i_3_n_0;
        release tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.sp_ram_i_i_4_n_0;
        release tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.wdata_i_IBUF;
        release tb.top_i.core_region_i.instr_mem.mem_gen_net.sp_ram_wrap_i.en_i_IBUF;
      `endif

    end
  endtask
`endif
